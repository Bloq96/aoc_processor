library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.GENERIC_FUNCTIONS.int2slv;
use work.GENERIC_FUNCTIONS.slv2int;

entity integer_divider is
    generic(
        DATA_LENGTH : natural);
    port(
        input_a : in std_logic_vector(11 downto 0);
        input_b : in std_logic_vector(9 downto 0);
        quotient : out std_logic_vector((DATA_LENGTH-1) downto 0);
        remainder : out std_logic_vector((DATA_LENGTH-1) downto 0));
end entity;

architecture behaviour_integer_division of integer_divider is
    constant MULTIPLIER_BITS : natural := (DATA_LENGTH - 12);    

    type division_lut_type is array((-512) to 511) of integer range
    (-(2**MULTIPLIER_BITS)) to (2**MULTIPLIER_BITS);
    constant DIV_LUT : division_lut_type := (
		-2048,-2052,-2056,-2060,-2064,-2068,-2072,-2076,
		-2081,-2085,-2089,-2093,-2097,-2101,-2106,-2110,
		-2114,-2118,-2123,-2127,-2131,-2136,-2140,-2144,
		-2149,-2153,-2158,-2162,-2166,-2171,-2175,-2180,
		-2185,-2189,-2194,-2198,-2203,-2208,-2212,-2217,
		-2222,-2226,-2231,-2236,-2241,-2245,-2250,-2255,
		-2260,-2265,-2270,-2275,-2280,-2284,-2289,-2294,
		-2300,-2305,-2310,-2315,-2320,-2325,-2330,-2335,
		-2341,-2346,-2351,-2356,-2362,-2367,-2372,-2378,
		-2383,-2389,-2394,-2399,-2405,-2411,-2416,-2422,
		-2427,-2433,-2439,-2444,-2450,-2456,-2461,-2467,
		-2473,-2479,-2485,-2491,-2497,-2503,-2509,-2515,
		-2521,-2527,-2533,-2539,-2545,-2551,-2558,-2564,
		-2570,-2576,-2583,-2589,-2595,-2602,-2608,-2615,
		-2621,-2628,-2635,-2641,-2648,-2655,-2661,-2668,
		-2675,-2682,-2689,-2696,-2703,-2709,-2717,-2724,
		-2731,-2738,-2745,-2752,-2759,-2767,-2774,-2781,
		-2789,-2796,-2804,-2811,-2819,-2826,-2834,-2842,
		-2849,-2857,-2865,-2873,-2881,-2889,-2897,-2905,
		-2913,-2921,-2929,-2937,-2945,-2954,-2962,-2970,
		-2979,-2987,-2996,-3005,-3013,-3022,-3031,-3039,
		-3048,-3057,-3066,-3075,-3084,-3093,-3102,-3112,
		-3121,-3130,-3139,-3149,-3158,-3168,-3178,-3187,
		-3197,-3207,-3216,-3226,-3236,-3246,-3256,-3267,
		-3277,-3287,-3297,-3308,-3318,-3329,-3339,-3350,
		-3361,-3372,-3383,-3393,-3404,-3416,-3427,-3438,
		-3449,-3461,-3472,-3484,-3495,-3507,-3519,-3531,
		-3542,-3554,-3567,-3579,-3591,-3603,-3616,-3628,
		-3641,-3654,-3666,-3679,-3692,-3705,-3718,-3732,
		-3745,-3758,-3772,-3785,-3799,-3813,-3827,-3841,
		-3855,-3869,-3884,-3898,-3913,-3927,-3942,-3957,
		-3972,-3987,-4002,-4018,-4033,-4049,-4064,-4080,
		-4096,-4112,-4128,-4145,-4161,-4178,-4194,-4211,
		-4228,-4245,-4263,-4280,-4297,-4315,-4333,-4351,
		-4369,-4387,-4406,-4424,-4443,-4462,-4481,-4500,
		-4520,-4539,-4559,-4579,-4599,-4619,-4640,-4660,
		-4681,-4702,-4723,-4745,-4766,-4788,-4810,-4832,
		-4855,-4877,-4900,-4923,-4946,-4970,-4993,-5017,
		-5041,-5066,-5090,-5115,-5140,-5165,-5191,-5217,
		-5243,-5269,-5296,-5323,-5350,-5377,-5405,-5433,
		-5461,-5490,-5519,-5548,-5578,-5607,-5638,-5668,
		-5699,-5730,-5761,-5793,-5825,-5858,-5891,-5924,
		-5958,-5992,-6026,-6061,-6096,-6132,-6168,-6205,
		-6242,-6279,-6317,-6355,-6394,-6433,-6473,-6513,
		-6554,-6595,-6637,-6679,-6722,-6765,-6809,-6853,
		-6899,-6944,-6991,-7037,-7085,-7133,-7182,-7232,
		-7282,-7333,-7384,-7437,-7490,-7544,-7598,-7654,
		-7710,-7767,-7825,-7884,-7944,-8004,-8066,-8128,
		-8192,-8257,-8322,-8389,-8456,-8525,-8595,-8666,
		-8738,-8812,-8886,-8962,-9039,-9118,-9198,-9279,
		-9362,-9447,-9533,-9620,-9709,-9800,-9892,-9986,
		-10082,-10180,-10280,-10382,-10486,-10592,-10700,-10810,
		-10923,-11038,-11155,-11275,-11398,-11523,-11651,-11782,
		-11916,-12053,-12193,-12336,-12483,-12633,-12788,-12945,
		-13107,-13273,-13443,-13618,-13797,-13981,-14170,-14364,
		-14564,-14769,-14980,-15197,-15420,-15650,-15888,-16132,
		-16384,-16644,-16913,-17190,-17476,-17772,-18079,-18396,
		-18725,-19065,-19418,-19784,-20165,-20560,-20972,-21400,
		-21845,-22310,-22795,-23302,-23831,-24385,-24966,-25575,
		-26214,-26887,-27594,-28340,-29127,-29959,-30840,-31775,
		-32768,-33825,-34953,-36158,-37449,-38836,-40330,-41943,
		-43691,-45590,-47663,-49932,-52429,-55188,-58254,-61681,
		-65536,-69905,-74898,-80660,-87381,-95325,-104858,-116508,
		-131072,-149797,-174763,-209715,-262144,-349525,-524288,-1048576,
		0,1048576,524288,349525,262144,209715,174763,149797,
		131072,116508,104858,95325,87381,80660,74898,69905,
		65536,61681,58254,55188,52429,49932,47663,45590,
		43691,41943,40330,38836,37449,36158,34953,33825,
		32768,31775,30840,29959,29127,28340,27594,26887,
		26214,25575,24966,24385,23831,23302,22795,22310,
		21845,21400,20972,20560,20165,19784,19418,19065,
		18725,18396,18079,17772,17476,17190,16913,16644,
		16384,16132,15888,15650,15420,15197,14980,14769,
		14564,14364,14170,13981,13797,13618,13443,13273,
		13107,12945,12788,12633,12483,12336,12193,12053,
		11916,11782,11651,11523,11398,11275,11155,11038,
		10923,10810,10700,10592,10486,10382,10280,10180,
		10082,9986,9892,9800,9709,9620,9533,9447,
		9362,9279,9198,9118,9039,8962,8886,8812,
		8738,8666,8595,8525,8456,8389,8322,8257,
		8192,8128,8066,8004,7944,7884,7825,7767,
		7710,7654,7598,7544,7490,7437,7384,7333,
		7282,7232,7182,7133,7085,7037,6991,6944,
		6899,6853,6809,6765,6722,6679,6637,6595,
		6554,6513,6473,6433,6394,6355,6317,6279,
		6242,6205,6168,6132,6096,6061,6026,5992,
		5958,5924,5891,5858,5825,5793,5761,5730,
		5699,5668,5638,5607,5578,5548,5519,5490,
		5461,5433,5405,5377,5350,5323,5296,5269,
		5243,5217,5191,5165,5140,5115,5090,5066,
		5041,5017,4993,4970,4946,4923,4900,4877,
		4855,4832,4810,4788,4766,4745,4723,4702,
		4681,4660,4640,4619,4599,4579,4559,4539,
		4520,4500,4481,4462,4443,4424,4406,4387,
		4369,4351,4333,4315,4297,4280,4263,4245,
		4228,4211,4194,4178,4161,4145,4128,4112,
		4096,4080,4064,4049,4033,4018,4002,3987,
		3972,3957,3942,3927,3913,3898,3884,3869,
		3855,3841,3827,3813,3799,3785,3772,3758,
		3745,3732,3718,3705,3692,3679,3666,3654,
		3641,3628,3616,3603,3591,3579,3567,3554,
		3542,3531,3519,3507,3495,3484,3472,3461,
		3449,3438,3427,3416,3404,3393,3383,3372,
		3361,3350,3339,3329,3318,3308,3297,3287,
		3277,3267,3256,3246,3236,3226,3216,3207,
		3197,3187,3178,3168,3158,3149,3139,3130,
		3121,3112,3102,3093,3084,3075,3066,3057,
		3048,3039,3031,3022,3013,3005,2996,2987,
		2979,2970,2962,2954,2945,2937,2929,2921,
		2913,2905,2897,2889,2881,2873,2865,2857,
		2849,2842,2834,2826,2819,2811,2804,2796,
		2789,2781,2774,2767,2759,2752,2745,2738,
		2731,2724,2717,2709,2703,2696,2689,2682,
		2675,2668,2661,2655,2648,2641,2635,2628,
		2621,2615,2608,2602,2595,2589,2583,2576,
		2570,2564,2558,2551,2545,2539,2533,2527,
		2521,2515,2509,2503,2497,2491,2485,2479,
		2473,2467,2461,2456,2450,2444,2439,2433,
		2427,2422,2416,2411,2405,2399,2394,2389,
		2383,2378,2372,2367,2362,2356,2351,2346,
		2341,2335,2330,2325,2320,2315,2310,2305,
		2300,2294,2289,2284,2280,2275,2270,2265,
		2260,2255,2250,2245,2241,2236,2231,2226,
		2222,2217,2212,2208,2203,2198,2194,2189,
		2185,2180,2175,2171,2166,2162,2158,2153,
		2149,2144,2140,2136,2131,2127,2123,2118,
		2114,2110,2106,2101,2097,2093,2089,2085,
		2081,2076,2072,2068,2064,2060,2056,2052);
    
    signal temp_a : integer := 0;
    signal temp_b : integer := 0;
    signal temp_q : integer := 0;
    signal temp_r : integer := 0;
    signal w_add_sub : std_logic;
    signal w_fix : std_logic;
    signal w_quot_fix : std_logic_vector((DATA_LENGTH-1) downto 0);
    signal w_quot_shft : std_logic_vector((DATA_LENGTH-1) downto
    0);
    signal w_rmdr_fix : std_logic_vector((DATA_LENGTH-1) downto 0);
    signal w_quot : std_logic_vector((DATA_LENGTH-1) downto 0);
    signal w_rmdr : std_logic_vector((DATA_LENGTH-1) downto 0);

    begin
        temp_a <= slv2int(input_a); 
        temp_b <= slv2int(input_b);
        w_quot_shft <= int2slv(temp_a*DIV_LUT(temp_b),DATA_LENGTH);
        w_quot((DATA_LENGTH-1) downto 12) <= (others
        => w_quot_shft(DATA_LENGTH-1));
        w_quot(11 downto 0) <= w_quot_shft((DATA_LENGTH-1) downto
        MULTIPLIER_BITS);
        temp_q <= slv2int(w_quot);
        temp_r <= temp_a-(temp_b*temp_q);
        w_rmdr <= int2slv(temp_r,DATA_LENGTH);
        quotient <= w_quot_fix when (w_fix = '1') else
                    w_quot;
        remainder <= w_rmdr_fix when (w_fix = '1') else
                     w_rmdr;
        w_add_sub <= '1' when ((input_b(9) xor w_rmdr(DATA_LENGTH-1))
        = '1') else
                 '0';
        w_quot_fix <= int2slv((temp_q-1),DATA_LENGTH) when 
                      (w_add_sub = '1') else
                      int2slv((temp_q+1),DATA_LENGTH);
        w_rmdr_fix <= int2slv((temp_r+temp_b),DATA_LENGTH) when 
                      (w_add_sub = '1') else
                      int2slv((temp_r-temp_b),DATA_LENGTH);
        w_fix <= '1' when ((abs(temp_r) >= abs(temp_b)) or
                 (((input_a(11) xor w_rmdr(DATA_LENGTH-1)) = '1') and
                 not(temp_r = 0))) else
                 '0';
end architecture;
